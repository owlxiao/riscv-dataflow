module Fetch
    import core_pkg::*;
(
    fetch_if.Fetch IO   ,
    CC_if.CoProcessor CC
);

endmodule
