module core
    import core_pkg::*;
(
    core_if.Master core_io
);

endmodule
