package core_pkg;
    import riscv_pkg::*;
endpackage
